paradicat@6/27
