tmtmmtm
