module demo(
	input  a,
	output b);
	
	assign b = ~a;
endmodule
