vvvvshs
dvjkds
